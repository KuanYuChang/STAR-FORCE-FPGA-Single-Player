module information_read_only (
input [16:0] addr,
output [11:0] pixel
);
parameter [11:0] mem [127999:0] = {
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hDDD,
12'h888,
12'h888,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h999,
12'h888,
12'h888,
12'h777,
12'h666,
12'h666,
12'h666,
12'h666,
12'h666,
12'h666,
12'h666,
12'h666,
12'h666,
12'h777,
12'h777,
12'h777,
12'h888,
12'h999,
12'hBBB,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hDDD,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'hDDD,
12'hEEE,
12'hDDD,
12'hEEE,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h888,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h888,
12'h999,
12'h999,
12'hAAA,
12'h999,
12'hAAA,
12'h555,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'h888,
12'h999,
12'hBBB,
12'hBBB,
12'hCCC,
12'hAAA,
12'h888,
12'h888,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'hAAA,
12'h444,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h666,
12'hCCC,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hEEE,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h999,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h111,
12'h000,
12'h333,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'hBBB,
12'hDDD,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hCCC,
12'h999,
12'h666,
12'h444,
12'h333,
12'h666,
12'h999,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h444,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'hCCC,
12'hCCC,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'hAAA,
12'h666,
12'h777,
12'h666,
12'h888,
12'h999,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hEEE,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h111,
12'h000,
12'h000,
12'h000,
12'h444,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h111,
12'h000,
12'h111,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hEEE,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hEEE,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h110,
12'hBBB,
12'hFFF,
12'hFFE,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'hDDD,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h111,
12'h111,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hEEE,
12'hFFF,
12'hFFF,
12'h444,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'hAAA,
12'hBBB,
12'hBBB,
12'hBBB,
12'hCCC,
12'hBBB,
12'hBBB,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h888,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hEED,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h888,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hDDD,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h666,
12'h666,
12'h666,
12'h888,
12'h888,
12'h888,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h888,
12'h888,
12'h777,
12'h777,
12'h888,
12'h888,
12'hBBB,
12'hEEE,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h111,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h111,
12'h333,
12'h222,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFE,
12'hEEE,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hCCC,
12'hBBB,
12'hDDD,
12'hDDD,
12'hEEE,
12'hDDD,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hDDD,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hBBB,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'hDDD,
12'hEEE,
12'hDDD,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hEEE,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'hCCC,
12'hDDD,
12'hCCC,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'hDDD,
12'hDDD,
12'hEEE,
12'hDDD,
12'hEEE,
12'hCCC,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h111,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFE,
12'hFFE,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hEEE,
12'hFFF,
12'hEEE,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFE,
12'hEEE,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h777,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'h888,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h888,
12'hFFF,
12'hDDD,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h554,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hCCC,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h666,
12'hFFF,
12'hEEE,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h999,
12'h666,
12'h555,
12'hAAA,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h999,
12'h777,
12'h777,
12'h777,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hDDD,
12'hCCC,
12'hBBB,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h111,
12'h777,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hCCC,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hCCC,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hBBB,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h999,
12'hBBB,
12'hCCC,
12'hBBB,
12'hBBB,
12'hAAA,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h777,
12'h888,
12'h999,
12'hBBB,
12'hAAA,
12'h888,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h777,
12'h888,
12'h999,
12'hAAA,
12'hAAA,
12'h999,
12'h999,
12'h888,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h333,
12'h444,
12'h444,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'hDDD,
12'hCCC,
12'hBBB,
12'hCCC,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDCD,
12'hDCD,
12'hCDD,
12'hCDD,
12'hCDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hDDD,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h011,
12'h000,
12'h101,
12'h000,
12'h112,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h110,
12'h000,
12'h222,
12'h000,
12'h000,
12'h111,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h551,
12'h995,
12'h220,
12'h000,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h555,
12'h999,
12'hAAA,
12'hBBB,
12'hAAA,
12'hAAA,
12'h888,
12'h444,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h333,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h000,
12'h000,
12'h000,
12'h444,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h555,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h444,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h444,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h110,
12'h110,
12'hDD6,
12'hEE8,
12'h995,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hEEE,
12'hFFF,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hDDD,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hDDD,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h101,
12'h000,
12'h000,
12'h100,
12'h551,
12'hFF6,
12'hEE4,
12'hFF8,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hEEE,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hAAA,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h999,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hAAA,
12'hDDD,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h999,
12'h000,
12'h888,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hAAA,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hAAA,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hBBB,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h100,
12'h000,
12'hCB6,
12'hFE4,
12'hEE2,
12'hFF5,
12'h771,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h111,
12'hCCC,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h333,
12'h999,
12'hFFF,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h666,
12'h666,
12'h666,
12'h777,
12'hBBB,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h888,
12'h555,
12'h666,
12'h777,
12'h777,
12'h999,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h666,
12'h777,
12'h888,
12'h777,
12'h777,
12'hAAA,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'hBBB,
12'h999,
12'h888,
12'h888,
12'h888,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h777,
12'h999,
12'h888,
12'h888,
12'h999,
12'hCCC,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h110,
12'h430,
12'hFF7,
12'hFE2,
12'hFF2,
12'hEE2,
12'hDD4,
12'h220,
12'h100,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hBBB,
12'hFFF,
12'hEEE,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hDDD,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hEEE,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h777,
12'hFFF,
12'h888,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h777,
12'hEEE,
12'hBBB,
12'h000,
12'h444,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h000,
12'h111,
12'h000,
12'h982,
12'hFE4,
12'hFE2,
12'hFF1,
12'hFF2,
12'hFF5,
12'h550,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'hDDD,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hCCC,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h220,
12'hEE5,
12'hFF3,
12'hFF2,
12'hFF2,
12'hFF2,
12'hEE2,
12'hCC5,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h112,
12'h000,
12'h100,
12'h652,
12'hFF6,
12'hEE3,
12'hCC1,
12'hEE3,
12'hEE1,
12'hFF3,
12'hEE6,
12'h440,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hEEE,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h100,
12'h210,
12'hBA6,
12'hEE7,
12'h891,
12'h550,
12'hBB3,
12'hFF4,
12'hDD1,
12'hFF5,
12'h992,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hEEE,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h011,
12'h000,
12'h000,
12'h100,
12'h320,
12'hFF8,
12'hEE8,
12'h010,
12'h000,
12'h550,
12'hFF5,
12'hFE3,
12'hFF4,
12'hEE5,
12'h220,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h121,
12'h000,
12'h210,
12'hBA3,
12'hFE5,
12'hEF7,
12'h9A4,
12'h000,
12'h110,
12'hEE6,
12'hFE4,
12'hFF3,
12'hFF5,
12'h772,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hBBB,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h888,
12'hEEE,
12'hFFF,
12'hDDD,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h555,
12'hDDD,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hEEE,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h122,
12'h000,
12'h000,
12'h320,
12'hFE5,
12'hEE3,
12'hFF7,
12'h340,
12'h120,
12'h000,
12'hA94,
12'hFE5,
12'hEE2,
12'hFF3,
12'hEF7,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hAAA,
12'hFFF,
12'hFFF,
12'h999,
12'h111,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h660,
12'hFF4,
12'hFF4,
12'hDD6,
12'h110,
12'h000,
12'h000,
12'h210,
12'hFF8,
12'hEE2,
12'hFF2,
12'hEE4,
12'h660,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'hEE6,
12'hFF3,
12'hEE2,
12'h880,
12'h440,
12'h330,
12'h440,
12'h220,
12'hBB3,
12'hFF3,
12'hFF1,
12'hFF3,
12'hDD4,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'h888,
12'h999,
12'hAAA,
12'hAAA,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h999,
12'h888,
12'hAAA,
12'hBBB,
12'hDDD,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h999,
12'hAAA,
12'h999,
12'hAAA,
12'hDDD,
12'hFFF,
12'hDDD,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBCC,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h113,
12'h000,
12'h550,
12'hFF5,
12'hEE2,
12'hFF2,
12'hFF4,
12'hEE4,
12'hEE4,
12'hFF5,
12'hFF4,
12'hEE2,
12'hFF1,
12'hFF1,
12'hEE0,
12'hFE4,
12'h440,
12'h010,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h112,
12'h110,
12'hBB3,
12'hDD2,
12'hEE2,
12'hFF3,
12'hFF5,
12'hFF5,
12'hFF4,
12'hFF5,
12'hFF5,
12'hFF4,
12'hEE1,
12'hFF1,
12'hFE1,
12'hFF3,
12'hBB5,
12'h110,
12'h000,
12'h001,
12'h001,
12'h000,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h111,
12'hEEE,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h221,
12'h330,
12'hEE5,
12'hFF4,
12'hFF6,
12'h770,
12'h430,
12'h651,
12'h550,
12'h430,
12'h551,
12'h440,
12'hAA1,
12'hFF4,
12'hFF2,
12'hEE2,
12'hFF6,
12'h440,
12'h000,
12'h001,
12'h000,
12'h011,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hEEE,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFE,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h882,
12'hFF5,
12'hDD3,
12'hFF8,
12'h110,
12'h000,
12'h000,
12'h000,
12'h110,
12'h000,
12'h110,
12'h430,
12'hFF6,
12'hED2,
12'hFF3,
12'hEE4,
12'h992,
12'h220,
12'h000,
12'h011,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h220,
12'hFF8,
12'hEE3,
12'hEF5,
12'h883,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h220,
12'hAA4,
12'hFF5,
12'hFF2,
12'hFE3,
12'hFE6,
12'h220,
12'h110,
12'h112,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h555,
12'hBBB,
12'hEEE,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hCCC,
12'hDDD,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h650,
12'hFE6,
12'hEE3,
12'hFF6,
12'h440,
12'h000,
12'h000,
12'h011,
12'h000,
12'h111,
12'h111,
12'h121,
12'h000,
12'h330,
12'hFF6,
12'hFF3,
12'hFF3,
12'hFF4,
12'h772,
12'h100,
12'h000,
12'h001,
12'h002,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'hCB3,
12'hFF4,
12'hFF4,
12'hCC4,
12'h000,
12'h010,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'hCC4,
12'hEE3,
12'hFF2,
12'hDD1,
12'hFF7,
12'h110,
12'h100,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h444,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h220,
12'hFF4,
12'hFE2,
12'hFF5,
12'h770,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h210,
12'h550,
12'hFF6,
12'hFE2,
12'hFF3,
12'hFF5,
12'h770,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h222,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hEEE,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h000,
12'h110,
12'h220,
12'hBB3,
12'hEE3,
12'hFF3,
12'hFE5,
12'h320,
12'h000,
12'h111,
12'h000,
12'h101,
12'h001,
12'h000,
12'h000,
12'h111,
12'h000,
12'h100,
12'h430,
12'hCC5,
12'hDD2,
12'hFF2,
12'hFF3,
12'hDD4,
12'h540,
12'h100,
12'h100,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h444,
12'h000,
12'h000,
12'h000,
12'h444,
12'h777,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h444,
12'h000,
12'h000,
12'h000,
12'h333,
12'h777,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h775,
12'h884,
12'hCC6,
12'hEE6,
12'hFF4,
12'hEE3,
12'hFF8,
12'h661,
12'h664,
12'h000,
12'h001,
12'h001,
12'h001,
12'h212,
12'h000,
12'h000,
12'h000,
12'h110,
12'h110,
12'hAA5,
12'hFF6,
12'hEE2,
12'hEF3,
12'hFE4,
12'hEE7,
12'hAA6,
12'h775,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h888,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hEEE,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h888,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hCCC,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hAAA,
12'h888,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h888,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBAB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h543,
12'hDDA,
12'hEE9,
12'hEE7,
12'hEF7,
12'hFF6,
12'hEE6,
12'hDE7,
12'hFFA,
12'hDDA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h111,
12'h000,
12'h110,
12'hEFB,
12'hDE6,
12'hEF6,
12'hEE4,
12'hFF7,
12'hED6,
12'hFF9,
12'hEEA,
12'hBB9,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hDDC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h221,
12'h552,
12'h773,
12'h560,
12'h550,
12'h550,
12'h550,
12'h661,
12'h562,
12'h220,
12'h332,
12'h000,
12'h111,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h121,
12'h110,
12'h230,
12'h551,
12'h560,
12'h660,
12'h660,
12'h761,
12'h661,
12'h552,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'h555,
12'h555,
12'h333,
12'h666,
12'h444,
12'h555,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h444,
12'h555,
12'h555,
12'h555,
12'h555,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h777,
12'h999,
12'h999,
12'hDDD,
12'hDDD,
12'hCCC,
12'hAAA,
12'h888,
12'h444,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'hDDD,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h666,
12'h555,
12'h444,
12'h444,
12'h444,
12'h444,
12'h555,
12'h555,
12'h555,
12'h555,
12'h777,
12'h777,
12'h777,
12'h888,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h444,
12'h555,
12'h444,
12'h444,
12'h444,
12'h444,
12'h555,
12'h555,
12'h555,
12'h666,
12'h555,
12'h777,
12'h666,
12'h666,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h555,
12'h555,
12'h555,
12'h444,
12'h444,
12'h555,
12'h555,
12'h555,
12'h666,
12'h666,
12'h666,
12'h666,
12'h777,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h555,
12'h555,
12'h555,
12'h444,
12'h444,
12'h555,
12'h555,
12'h666,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h443,
12'h666,
12'h554,
12'h444,
12'h444,
12'h555,
12'h555,
12'h555,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h100,
12'h000,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h010,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h010,
12'h010,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h101,
12'h001,
12'h102,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h111,
12'h000,
12'h000,
12'h011,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hDDC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h011,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h777,
12'hCCC,
12'hDDD,
12'hCCC,
12'hBBB,
12'hDDD,
12'hCCC,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCC,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hDDD,
12'hDDD,
12'hDDD,
12'hCDD,
12'hCDD,
12'hCDD,
12'hCDD,
12'hDDD,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCC,
12'hCCC,
12'hCCD,
12'hCCD,
12'hDDD,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hBBB,
12'hCCC,
12'hDDD,
12'hCCD,
12'hCCC,
12'hDDD,
12'hDDD,
12'hDCD,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCC,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCD,
12'hDCD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCDD,
12'hCDD,
12'hCDD,
12'hCDC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hEEE,
12'h888,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'h555,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h010,
12'h000,
12'h442,
12'h441,
12'h440,
12'h440,
12'h320,
12'h430,
12'h330,
12'h440,
12'h450,
12'h340,
12'h551,
12'h441,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h777,
12'h888,
12'hAAA,
12'hBBB,
12'h999,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h666,
12'h999,
12'hBBB,
12'hBBB,
12'hBBB,
12'hAAA,
12'h999,
12'h666,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'h888,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h555,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEED,
12'hEFD,
12'hEFA,
12'hEE8,
12'hFE8,
12'hFE8,
12'hFF9,
12'hFF9,
12'hDE7,
12'hFF9,
12'hEF9,
12'hEF9,
12'hEE8,
12'hEE9,
12'hFFA,
12'hFFA,
12'hDD8,
12'hBA6,
12'h652,
12'h330,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'hCCC,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hDDD,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h998,
12'h997,
12'hDD8,
12'hDD6,
12'hFF5,
12'hFF5,
12'hDD5,
12'hEE7,
12'hFF9,
12'hDD7,
12'hFF9,
12'hEF8,
12'hEE7,
12'hEE6,
12'hEF7,
12'hFF7,
12'hEF6,
12'hEE5,
12'hFF6,
12'hFE6,
12'hDC5,
12'h550,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hCCC,
12'hBBB,
12'h000,
12'h555,
12'hAAA,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h444,
12'h999,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h999,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hBBB,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h999,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h888,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h450,
12'hFF7,
12'hFF4,
12'hEE3,
12'hFF6,
12'h660,
12'h551,
12'h440,
12'h330,
12'h561,
12'h771,
12'h881,
12'hAA3,
12'hDE6,
12'hFF7,
12'hEE5,
12'hED3,
12'hFF4,
12'hFF4,
12'hFF6,
12'hCC7,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hCCC,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h777,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hEEE,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h666,
12'h666,
12'h666,
12'h777,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hEEE,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h333,
12'h777,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hEEE,
12'hFFF,
12'hBBB,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hCCC,
12'hAAA,
12'h999,
12'h999,
12'h999,
12'h777,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h888,
12'h888,
12'h999,
12'h999,
12'hBBB,
12'hCCC,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h440,
12'hFF7,
12'hEE3,
12'hEE3,
12'hFE7,
12'h110,
12'h000,
12'h000,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h010,
12'h551,
12'hBB5,
12'hFF7,
12'hFE4,
12'hEE3,
12'hEE3,
12'hFF6,
12'hEE8,
12'h220,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hBCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hEEE,
12'hBBB,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h450,
12'hDD5,
12'hEE3,
12'hFF5,
12'hEE8,
12'h330,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h650,
12'hFF8,
12'hFF6,
12'hFF4,
12'hDE3,
12'hFF5,
12'hED8,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hEEE,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h450,
12'hEF7,
12'hFF4,
12'hEE4,
12'hFE8,
12'h430,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEE9,
12'hFF7,
12'hFF3,
12'hEE2,
12'hFF6,
12'hDC6,
12'h210,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hCDC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h440,
12'hFF7,
12'hFE4,
12'hFE5,
12'hFE9,
12'h100,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h000,
12'h112,
12'h000,
12'h000,
12'hEE8,
12'hDD2,
12'hFF2,
12'hED2,
12'hFE6,
12'h551,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hEEE,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h555,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hCCC,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h440,
12'hFF7,
12'hEE4,
12'hEE4,
12'hEE9,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h330,
12'hFF6,
12'hEE2,
12'hFF2,
12'hEE4,
12'hDD7,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hDDD,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h340,
12'hFF7,
12'hEE4,
12'hFE5,
12'hFE9,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'hCC4,
12'hEE4,
12'hFF2,
12'hEE2,
12'hEE7,
12'h330,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hEEE,
12'hFFF,
12'hDDD,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h330,
12'hFF7,
12'hFE3,
12'hFE5,
12'hFE9,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h661,
12'hEE6,
12'hFF3,
12'hFF3,
12'hFF6,
12'h772,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hEEE,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hEEE,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h777,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h330,
12'hFF7,
12'hFE3,
12'hFE4,
12'hFE9,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'hEE8,
12'hFE4,
12'hFF3,
12'hFF4,
12'h9A3,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hEEE,
12'hFFF,
12'hDDD,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h330,
12'hFF7,
12'hFE3,
12'hFE4,
12'hFE9,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDD8,
12'hFF4,
12'hEE2,
12'hFF4,
12'hBB3,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hEEE,
12'h111,
12'h111,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hEEE,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'h888,
12'h888,
12'h777,
12'h777,
12'h777,
12'h888,
12'h888,
12'h999,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h330,
12'hFF7,
12'hFE3,
12'hFE4,
12'hFE9,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'hCC7,
12'hFF5,
12'hEE2,
12'hFF5,
12'hAA3,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hAAA,
12'hEEE,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hEEE,
12'hCCC,
12'h777,
12'h999,
12'hBBB,
12'hAAA,
12'hCCC,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hDDD,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hEEE,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h330,
12'hFF7,
12'hFE3,
12'hFE3,
12'hFE8,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'hDC7,
12'hFF5,
12'hFE3,
12'hFF6,
12'h982,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h330,
12'hFF7,
12'hFF3,
12'hFE3,
12'hFE8,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFE8,
12'hFE4,
12'hEE3,
12'hEE6,
12'h762,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h222,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h888,
12'h888,
12'h888,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h330,
12'hEE6,
12'hFF4,
12'hFE3,
12'hEE8,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h100,
12'hFE7,
12'hFF4,
12'hEE3,
12'hFE9,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h330,
12'hEE7,
12'hFE3,
12'hFF4,
12'hFF8,
12'h210,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h772,
12'hFE6,
12'hEE3,
12'hFF5,
12'hBA6,
12'h100,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h555,
12'h000,
12'hBBB,
12'hEEE,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h444,
12'hFFF,
12'hDDD,
12'hEEE,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hEEE,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h330,
12'hFF7,
12'hEE3,
12'hEE3,
12'hFF7,
12'h330,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEE7,
12'hFF5,
12'hEE4,
12'hFF7,
12'h441,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'hCCC,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h440,
12'hFF7,
12'hFF3,
12'hFE3,
12'hEE6,
12'h430,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h772,
12'hFF6,
12'hDD3,
12'hEE6,
12'hBA4,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'hDDD,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hDDD,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hEEE,
12'hEEE,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h440,
12'hFE6,
12'hFE3,
12'hFF3,
12'hEE6,
12'h430,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h440,
12'hFF7,
12'hFF6,
12'hDE5,
12'hFF9,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'h999,
12'h000,
12'h111,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h550,
12'hFF6,
12'hEE2,
12'hEE2,
12'hFF5,
12'h770,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'hAA5,
12'hFF8,
12'hDE5,
12'hEE5,
12'hFF8,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hEEE,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h771,
12'hFF6,
12'hFE2,
12'hFE1,
12'hFF5,
12'hBB3,
12'h440,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h220,
12'h662,
12'h9A4,
12'hEF8,
12'hDE6,
12'hFF7,
12'hEE7,
12'hEE9,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hEEE,
12'hFFF,
12'hEEE,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h555,
12'h111,
12'h000,
12'h000,
12'h444,
12'h555,
12'hCCC,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hDDD,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h664,
12'hCC6,
12'hEE5,
12'hFE3,
12'hFF3,
12'hEE4,
12'hFF7,
12'hFF9,
12'hEEA,
12'hEEA,
12'hCC9,
12'hCC8,
12'hDC9,
12'hEEA,
12'hEE9,
12'hEE9,
12'hEE8,
12'hEF8,
12'hFF8,
12'hDD6,
12'h994,
12'h100,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h555,
12'h999,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h999,
12'h888,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hCCC,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h666,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h777,
12'h444,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hDDD,
12'hAAA,
12'h777,
12'h555,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hBBB,
12'h888,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h777,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h999,
12'h888,
12'h666,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h666,
12'hAAA,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h888,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h000,
12'h000,
12'hBBB,
12'hEEC,
12'hFEA,
12'hFE8,
12'hFE6,
12'hFE6,
12'hEE6,
12'hEE6,
12'hEE7,
12'hFF8,
12'hFE8,
12'hEF7,
12'hEE7,
12'hEE7,
12'hFF8,
12'hFF9,
12'hFFA,
12'hEEA,
12'hCC9,
12'h664,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h998,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h889,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h554,
12'h552,
12'h551,
12'h550,
12'h660,
12'h661,
12'h771,
12'h882,
12'h983,
12'h882,
12'h9A3,
12'hAA3,
12'hAA3,
12'h993,
12'h762,
12'h330,
12'h100,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h555,
12'h555,
12'h555,
12'h555,
12'h333,
12'h666,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h444,
12'h444,
12'h555,
12'h555,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h666,
12'h999,
12'hDDD,
12'hEEE,
12'hCCC,
12'hCCC,
12'hBBB,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h999,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'h555,
12'h444,
12'h444,
12'h444,
12'h444,
12'h555,
12'h555,
12'h666,
12'h666,
12'h666,
12'h777,
12'h777,
12'h777,
12'h444,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h555,
12'h555,
12'h444,
12'h444,
12'h444,
12'h555,
12'h666,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h666,
12'h666,
12'h555,
12'h666,
12'h555,
12'h666,
12'h555,
12'h444,
12'h444,
12'h444,
12'h555,
12'h555,
12'h555,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h777,
12'h999,
12'hBBB,
12'hCCC,
12'hDDD,
12'hDDD,
12'hCCC,
12'hAAA,
12'h666,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h555,
12'h444,
12'h444,
12'h444,
12'h555,
12'h333,
12'h666,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h555,
12'h444,
12'h555,
12'h444,
12'h555,
12'h555,
12'h555,
12'h555,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h555,
12'h555,
12'h555,
12'h444,
12'h444,
12'h777,
12'h444,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h887,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hDDD,
12'hDDD,
12'hCCC,
12'hBBB,
12'hDDD,
12'hDDD,
12'hDDD,
12'hCCC,
12'hDDD,
12'hCCC,
12'hCCC,
12'hEEE,
12'hCCC,
12'hCCC,
12'hCCC,
12'hDCD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hCCC,
12'hCCC,
12'hDDD,
12'hDDD,
12'hCCD,
12'hCCC,
12'hCCD,
12'hDCD,
12'hDDD,
12'hDDD,
12'hCCC,
12'hCCC,
12'hCCC,
12'hDDD,
12'hDDD,
12'hDDD,
12'hCCC,
12'hCCC,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDC,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hABA,
12'hBBB,
12'hEEE,
12'hBBC,
12'hCCC,
12'hDDE,
12'hCCD,
12'hDDE,
12'hDDD,
12'hCCC,
12'hCCC,
12'hDDD,
12'hDDD,
12'hDDD,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hDDD,
12'hCCC,
12'hCCC,
12'hDDD,
12'hCCC,
12'hEEE,
12'hCCC,
12'hCCC,
12'hCCC,
12'hDDD,
12'hCCC,
12'hDDE,
12'hCCD,
12'hDCD,
12'hDDD,
12'hDCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hCCC,
12'hDDC,
12'hDDC,
12'hDDD,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h221,
12'h010,
12'h220,
12'h110,
12'h220,
12'h120,
12'h000,
12'h110,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h220,
12'h110,
12'h220,
12'h110,
12'h110,
12'h220,
12'h110,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDC,
12'h110,
12'h110,
12'h452,
12'h996,
12'h995,
12'h994,
12'h883,
12'h883,
12'h883,
12'h894,
12'hAA7,
12'h885,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h776,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h664,
12'h996,
12'h995,
12'h883,
12'h883,
12'h894,
12'hAA6,
12'h886,
12'h443,
12'h110,
12'h110,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'hCCC,
12'hAAA,
12'h999,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h999,
12'h888,
12'h888,
12'hCCC,
12'hDDD,
12'h555,
12'h000,
12'h444,
12'hFFF,
12'hDDD,
12'hBBB,
12'h999,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h999,
12'h888,
12'hAAA,
12'hBBB,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hAAA,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hDDD,
12'hAAA,
12'h777,
12'h333,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h999,
12'hAAA,
12'h999,
12'h888,
12'h888,
12'h999,
12'hAAA,
12'h999,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'h999,
12'h999,
12'h888,
12'h999,
12'h999,
12'hAAA,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCB,
12'h010,
12'h221,
12'hBB9,
12'hEEA,
12'hEF9,
12'hFE7,
12'hFF6,
12'hFE4,
12'hFF5,
12'hFF6,
12'hEE8,
12'hEFB,
12'h775,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h220,
12'hED9,
12'hFEA,
12'h540,
12'h331,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFC,
12'hDD9,
12'hFE8,
12'hEE5,
12'hFF6,
12'hEE6,
12'hFF8,
12'hFEA,
12'hCB9,
12'h221,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hEEE,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hAAA,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCDC,
12'h110,
12'h010,
12'h231,
12'h440,
12'h660,
12'hDD5,
12'hFF5,
12'hFE2,
12'hFF3,
12'hEE4,
12'h881,
12'h450,
12'h010,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h330,
12'h661,
12'hFE8,
12'hFE7,
12'hCC6,
12'h220,
12'h000,
12'h000,
12'h000,
12'h100,
12'h000,
12'h000,
12'h000,
12'h000,
12'h330,
12'h440,
12'hEE6,
12'hFF4,
12'hFE4,
12'hFF6,
12'h881,
12'h440,
12'h220,
12'h000,
12'h111,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h667,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hAAA,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFE,
12'hDDC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hCCC,
12'hBBB,
12'h999,
12'h888,
12'h999,
12'hAAA,
12'hCCC,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h444,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDED,
12'h010,
12'h000,
12'h000,
12'h110,
12'h210,
12'h660,
12'hFF6,
12'hFE3,
12'hFF3,
12'hFF4,
12'h881,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'hAA3,
12'hFF6,
12'hEE4,
12'hFF6,
12'h330,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h320,
12'hEE6,
12'hFE5,
12'hEE5,
12'hAA4,
12'h330,
12'h110,
12'h110,
12'h111,
12'h001,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hEEE,
12'h666,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h888,
12'hFFF,
12'hDDD,
12'h888,
12'h333,
12'hFFF,
12'hFFF,
12'h777,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h555,
12'hAAA,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h333,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEED,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h110,
12'hED7,
12'hFE4,
12'hFF3,
12'hFF4,
12'hCC4,
12'h220,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h320,
12'hFF7,
12'hFF4,
12'hFF3,
12'hEF4,
12'h994,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h540,
12'hFF7,
12'hEE4,
12'hFF6,
12'h440,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'h888,
12'h444,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hEEE,
12'hEEE,
12'hFFF,
12'hEEE,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDED,
12'h010,
12'h000,
12'h000,
12'h000,
12'h000,
12'h210,
12'h993,
12'hEE4,
12'hFE2,
12'hFF3,
12'hEE5,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h222,
12'h000,
12'h110,
12'hA94,
12'hFF6,
12'hDD1,
12'hFF1,
12'hFF4,
12'hEE7,
12'h320,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h992,
12'hFF6,
12'hFF5,
12'hDD5,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hEEF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h430,
12'hFF6,
12'hEE2,
12'hFF2,
12'hFF5,
12'h661,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h220,
12'hFE8,
12'hED4,
12'hFF3,
12'hEE0,
12'hFF3,
12'hFF6,
12'h761,
12'h210,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h220,
12'hFE7,
12'hEE5,
12'hFF6,
12'h660,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFE,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hEEE,
12'hFFF,
12'h888,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h220,
12'hDD5,
12'hFE3,
12'hEE1,
12'hFE4,
12'hBB5,
12'h110,
12'h110,
12'h110,
12'h000,
12'h000,
12'h000,
12'h110,
12'h771,
12'hFF7,
12'hFE5,
12'hFF4,
12'hFF3,
12'hFF2,
12'hFF4,
12'hCC4,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h540,
12'hFE6,
12'hED4,
12'hFE7,
12'h330,
12'h220,
12'h000,
12'h000,
12'h000,
12'h001,
12'h101,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'h334,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h881,
12'hFF5,
12'hFE2,
12'hEE3,
12'hFF8,
12'h220,
12'h000,
12'h221,
12'h010,
12'h000,
12'h000,
12'h110,
12'hDD6,
12'hEE6,
12'hFE7,
12'h770,
12'hFE4,
12'hEE2,
12'hFF3,
12'hEE5,
12'h330,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'hA94,
12'hED4,
12'hFE6,
12'hBA5,
12'h110,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h887,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hEEE,
12'hCCC,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h440,
12'hFF7,
12'hFF4,
12'hFE3,
12'hFF6,
12'h550,
12'h000,
12'h111,
12'h000,
12'h010,
12'h000,
12'h440,
12'hFF7,
12'hEE6,
12'hDD8,
12'h210,
12'hCC3,
12'hFF4,
12'hEE2,
12'hFF5,
12'h994,
12'h110,
12'h110,
12'h100,
12'h000,
12'h000,
12'h220,
12'hEE7,
12'hFE5,
12'hFE6,
12'h440,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h888,
12'hFFF,
12'hFFE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h220,
12'hDC6,
12'hFE4,
12'hFF3,
12'hFF5,
12'hAA3,
12'h000,
12'h000,
12'h000,
12'h000,
12'h120,
12'hAB5,
12'hFF7,
12'hFF7,
12'h652,
12'h110,
12'h771,
12'hFF6,
12'hEE2,
12'hFF5,
12'hDD7,
12'h220,
12'h110,
12'h000,
12'h000,
12'h000,
12'h450,
12'hFF7,
12'hFE6,
12'hFE7,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h222,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h883,
12'hFE4,
12'hFF3,
12'hFF3,
12'hEE5,
12'h110,
12'h000,
12'h000,
12'h000,
12'h230,
12'hEF8,
12'hFE6,
12'hFE7,
12'h110,
12'h010,
12'h320,
12'hEE6,
12'hFF4,
12'hEF3,
12'hFF6,
12'h660,
12'h110,
12'h000,
12'h000,
12'h110,
12'hAB4,
12'hFF6,
12'hEE6,
12'hAA4,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEED,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h100,
12'h430,
12'hEE5,
12'hFF2,
12'hFF2,
12'hFF5,
12'h440,
12'h110,
12'h000,
12'h110,
12'h893,
12'hFF7,
12'hFF7,
12'h882,
12'h220,
12'h000,
12'h000,
12'hAA4,
12'hFF5,
12'hEE2,
12'hFF4,
12'hCC4,
12'h000,
12'h000,
12'h000,
12'h230,
12'hEF6,
12'hEE5,
12'hEE7,
12'h440,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'hCC4,
12'hFF4,
12'hEE2,
12'hFF4,
12'h984,
12'h100,
12'h000,
12'h220,
12'hEE7,
12'hEE6,
12'hFF9,
12'h330,
12'h110,
12'h000,
12'h000,
12'h440,
12'hEE5,
12'hFF3,
12'hFF2,
12'hFF5,
12'h210,
12'h000,
12'h000,
12'h551,
12'hEE5,
12'hEE5,
12'hDD7,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h888,
12'hAAA,
12'h888,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h999,
12'h999,
12'h999,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h210,
12'h882,
12'hFF6,
12'hFE2,
12'hFE4,
12'hDD7,
12'h220,
12'h000,
12'h662,
12'hFE6,
12'hEE6,
12'hBB6,
12'h210,
12'h000,
12'h000,
12'h000,
12'h120,
12'hCC4,
12'hFF4,
12'hFE2,
12'hFF4,
12'h994,
12'h110,
12'h110,
12'hBA5,
12'hEF5,
12'hFF6,
12'h773,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h220,
12'h440,
12'hEE6,
12'hFE4,
12'hFE4,
12'hFE7,
12'h440,
12'h110,
12'hCC6,
12'hFE6,
12'hFF7,
12'h441,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h771,
12'hFE6,
12'hFE3,
12'hFE4,
12'hFF8,
12'h330,
12'h330,
12'hFF9,
12'hFF7,
12'hED6,
12'h220,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hEEE,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEED,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h221,
12'h210,
12'hCC6,
12'hFF5,
12'hFE3,
12'hFF6,
12'h770,
12'h450,
12'hFF8,
12'hEE5,
12'hDC5,
12'h110,
12'h110,
12'h001,
12'h000,
12'h000,
12'h000,
12'h220,
12'hFE7,
12'hFE4,
12'hFE3,
12'hFE6,
12'h550,
12'h660,
12'hFE8,
12'hED6,
12'hCB5,
12'h220,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h333,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h100,
12'h873,
12'hFE5,
12'hFF2,
12'hFF3,
12'hCC1,
12'hBA0,
12'hFF6,
12'hFF7,
12'h660,
12'h220,
12'h000,
12'h000,
12'h001,
12'h001,
12'h000,
12'h220,
12'h993,
12'hFF4,
12'hFE2,
12'hEE3,
12'hDC2,
12'hAA0,
12'hFE6,
12'hFF7,
12'h661,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h100,
12'h430,
12'hFF6,
12'hEF2,
12'hFE1,
12'hFF2,
12'hEE2,
12'hFF5,
12'hDD7,
12'h330,
12'h210,
12'h110,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h440,
12'hFF6,
12'hFF3,
12'hFE2,
12'hEE1,
12'hFF3,
12'hFF5,
12'hDD7,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'hDD5,
12'hFF4,
12'hFE1,
12'hFF2,
12'hEE2,
12'hFF5,
12'h983,
12'h110,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'hCC4,
12'hFF4,
12'hFF2,
12'hFE1,
12'hEE1,
12'hEE4,
12'hAA4,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFE,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h777,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h222,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h100,
12'h000,
12'h220,
12'h872,
12'hFF6,
12'hEE2,
12'hFF1,
12'hEF3,
12'hFF6,
12'h330,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h220,
12'h661,
12'hFF6,
12'hEE2,
12'hFF2,
12'hDD0,
12'hFF6,
12'h440,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hEEE,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hEEE,
12'hEEE,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h321,
12'h330,
12'hFE7,
12'hFE3,
12'hEE2,
12'hFF5,
12'hBB4,
12'h110,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h220,
12'hEE8,
12'hDE2,
12'hFF2,
12'hFF3,
12'hDE5,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h110,
12'hCC7,
12'hFE5,
12'hEE4,
12'hFF6,
12'h440,
12'h220,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h220,
12'h994,
12'hFF6,
12'hDD2,
12'hFF6,
12'h771,
12'h220,
12'h111,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hEEE,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h555,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hBBB,
12'h777,
12'h777,
12'h777,
12'h777,
12'h999,
12'hCCC,
12'hFFE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h763,
12'hEE6,
12'hFF6,
12'hBC6,
12'h120,
12'h111,
12'h000,
12'h000,
12'h110,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h330,
12'hFF7,
12'hEE6,
12'hEE8,
12'h220,
12'h220,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h111,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h888,
12'hEEE,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'hFFE,
12'hFFF,
12'hDDD,
12'h444,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h110,
12'hFF9,
12'hEE8,
12'h551,
12'h120,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'hAB5,
12'hFF9,
12'hA96,
12'h100,
12'h221,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hEED,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h333,
12'hAAA,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h442,
12'h110,
12'h000,
12'h011,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h110,
12'h653,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h333,
12'h666,
12'h666,
12'h666,
12'h776,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h221,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hCCC,
12'hDDD,
12'hBBB,
12'hBCC,
12'hCDD,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCC,
12'hCCC,
12'hCCC,
12'hDDD,
12'hCCC,
12'hDDD,
12'hCDD,
12'hCCC,
12'hDCC,
12'hDCC,
12'hDCC,
12'hDDC,
12'hDDD,
12'hCDD,
12'hCDD,
12'hCDD,
12'hDDC,
12'hDDC,
12'hDDC,
12'hCCD,
12'hCCD,
12'hCCD,
12'hCCC,
12'hDDD,
12'hCCC,
12'hDCD,
12'hCCD,
12'hDDD,
12'hDDD,
12'hDDC,
12'hDDC,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'hDDD,
12'h222,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h001,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h333,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hDDD,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h777,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'hBBB,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h555,
12'h999,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hEEE,
12'hEEE,
12'hEEE,
12'hEEE,
12'hDDD,
12'hEEE,
12'hFFF,
12'h444,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'hBBB,
12'h665,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h555,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hBBB,
12'h999,
12'hBBB,
12'hDDD,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'hFFF,
12'hFFF,
12'hDDD,
12'h999,
12'h000,
12'h333,
12'h777,
12'hDDD,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h888,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hEEE,
12'h999,
12'h000,
12'h111,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'h333,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hBBB,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hEEE,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hEEE,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hEEE,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hEEE,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hDDD,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hEEE,
12'hFFF,
12'h999,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h777,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hEEE,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hEEE,
12'h555,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'h999,
12'h111,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hEEE,
12'h444,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'h444,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h222,
12'h555,
12'h333,
12'h999,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hEEE,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h333,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hBBB,
12'hDDD,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'hCCC,
12'hCCC,
12'hEEE,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hAAA,
12'hBBB,
12'hBBB,
12'hBBB,
12'hFFF,
12'hFFF,
12'h666,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hAAA,
12'hAAA,
12'hCCC,
12'h888,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hEEE,
12'hFFF,
12'h888,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h999,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'hCCC,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'h555,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h555,
12'hEEE,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hDDD,
12'hFFF,
12'h333,
12'hFFF,
12'hFFF,
12'h444,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'hFFF,
12'h999,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h999,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hFFF,
12'hFFF,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hEEE,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hEEE,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hEEE,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h444,
12'hFFF,
12'hEEE,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h555,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hAAA,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hDDD,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hBBB,
12'h333,
12'h111,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'hFFF,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hEEE,
12'hFFF,
12'hBBB,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hEEE,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'hFFF,
12'hFFF,
12'hFFF,
12'h888,
12'h777,
12'h555,
12'h666,
12'hAAA,
12'hFFF,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hEEE,
12'h333,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h666,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hEEE,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hCCC,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h777,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h555,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hCCC,
12'h000,
12'h000,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hEEE,
12'hFFF,
12'hFFF,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hEEE,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h444,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h222,
12'h888,
12'h888,
12'h777,
12'h777,
12'h999,
12'h888,
12'h888,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hCCC,
12'hDDD,
12'hDDD,
12'hEEE,
12'hDDD,
12'h999,
12'h555,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hBBB,
12'hAAA,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h777,
12'hDDD,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'h888,
12'hAAA,
12'h999,
12'h999,
12'h000,
12'h111,
12'h000,
12'h777,
12'h777,
12'h888,
12'h888,
12'h777,
12'h888,
12'h888,
12'h444,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h111,
12'h555,
12'h888,
12'h777,
12'h777,
12'h888,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h111,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000
};
assign pixel = mem[addr];
endmodule
